`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Caite Sklar
// 
// Module Name: alu_tb
// Project Name: CPU-Core
// Target Devices: 
// Tool Versions: 
// Description: Tests all 7 alu operations.
// 
// Dependencies: alu
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module alu_tb;
    reg [15:0] a;
    reg [15:0] b;
    reg [3:0] sel;
    wire [15:0] out;
    
    alu alu (
        .in0(a),
        .in1(b),
        .select(sel),
        .out(out)
    );

    initial begin
        a = 13;
        b = 6;
        
        sel = 0;
        #2 assert(out == a) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 1;
        #2 assert(out == b) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 2;
        #2 assert(out == (a + b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 3;
        #2 assert(out == (a - b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);
        
        #5 sel = 4;
        #2 assert(out == (a * b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 5;
        #2 assert(out == (a / b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 6;
        #2 assert(out == (a & b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 7;
        #2 assert(out == (a | b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 8;
        #2 assert(out == (a ^ b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 9;
        #2 assert(out == (a << b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 10;
        #2 assert(out == (a >> b)) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);

        #5 sel = 11;
        #2 assert(out == 0) else $fatal(1, "Unexpected result: sel=%b a=%b b=%b out=%b", sel, a, b, out);
  
        #5;
         // No fatal errors
        $display ("*** ALU Testbench Passed");
        $finish;
    end

endmodule